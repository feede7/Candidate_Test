------------------------------------------------------------------------------
-- Company: Satellogic S.A
--
-- File: axi_spi.vhdl
-- Description: 
--
-- AXI-SPI device for new candidates
--
-- Author: Andres Demski
--
--------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;


entity axi_spi  is
    generic (
        C_AXI_DATA_WIDTH : integer :=32;
        C_AXI_ADDR_WIDTH : integer :=4
    );
    port (
        -- AXI4-Lite Slave Port
        AXI_ACLK             : in std_logic;
        AXI_ARESETN          : in std_logic;
        AXI_AWADDR           : in std_logic_vector(C_AXI_ADDR_WIDTH-1 downto 0);
        AXI_AWVALID          : in std_logic;
        AXI_AWREADY          : out std_logic;
        AXI_WDATA            : in std_logic_vector(C_AXI_DATA_WIDTH-1 downto 0);
        AXI_WSTRB            : in std_logic_vector(C_AXI_DATA_WIDTH/8-1 downto 0);           
        AXI_WVALID           : in std_logic;
        AXI_WREADY           : out std_logic;
        AXI_BRESP            : out std_logic_vector(1 downto 0);
        AXI_BVALID           : out std_logic;
        AXI_BREADY           : in std_logic;
        AXI_ARADDR           : in std_logic_vector(C_AXI_ADDR_WIDTH-1 downto 0);
        AXI_ARVALID          : in std_logic;
        AXI_ARREADY          : out std_logic;
        AXI_RDATA            : out std_logic_vector(C_AXI_DATA_WIDTH-1 downto 0);
        AXI_RRESP            : out std_logic_vector(1 downto 0);
        AXI_RVALID           : out std_logic;
        AXI_RREADY           : in std_logic;

        -- SPI Signals
        MOSI                 : out std_logic;
        MISO                 : in std_logic;
        SCLK                 : out std_logic;
        CSn                  : out std_logic;
        INT                  : out std_logic
    );
end axi_spi;

architecture arch_imp of axi_spi is

    signal WDATA  	: std_logic_vector(C_AXI_DATA_WIDTH-1 downto 0);
    signal RDATA  	: std_logic_vector(C_AXI_DATA_WIDTH-1 downto 0);
    signal RADDR  	: std_logic_vector(C_AXI_ADDR_WIDTH -1 downto 0);
    signal WADDR  	: std_logic_vector(C_AXI_ADDR_WIDTH -1 downto 0);
    signal WENA   	: std_logic;                           
    signal RENA   	: std_logic;
begin

    AXI_REGISTERS: entity work.axi_lite_slave_int
        generic map(
            C_S_AXI_DATA_WIDTH     => C_AXI_DATA_WIDTH,
            C_S_AXI_ADDR_WIDTH     => C_AXI_ADDR_WIDTH)
        port map (
            WDATA_O                => WDATA,
            RDATA_I                => RDATA,
            WENA_O                 => WENA,
            RENA_O                 => RENA,
            RADDR_O                => RADDR,
            WADDR_O                => WADDR,
            S_AXI_ACLK             => AXI_ACLK,
            S_AXI_ARESETN          => AXI_ARESETN,
            S_AXI_AWADDR           => AXI_AWADDR,
            S_AXI_AWVALID          => AXI_AWVALID,
            S_AXI_AWREADY          => AXI_AWREADY,
            S_AXI_WDATA            => AXI_WDATA,
            S_AXI_WSTRB            => AXI_WSTRB,
            S_AXI_WVALID           => AXI_WVALID,
            S_AXI_WREADY           => AXI_WREADY,
            S_AXI_BRESP            => AXI_BRESP,
            S_AXI_BVALID           => AXI_BVALID,
            S_AXI_BREADY           => AXI_BREADY,
            S_AXI_ARADDR           => AXI_ARADDR,
            S_AXI_ARVALID          => AXI_ARVALID,
            S_AXI_ARREADY          => AXI_ARREADY,
            S_AXI_RDATA            => AXI_RDATA,
            S_AXI_RRESP            => AXI_RRESP,
            S_AXI_RVALID           => AXI_RVALID,
            S_AXI_RREADY           => AXI_RREADY
        );    

    ---------------------------------------------------------
    -- Intanciar CORE AQUI!
    
	--    +-----+                                             +-----+
	--    |     |                                             |     |
	--    |     |      +----------------------------+         |     |
	--    |     |      |       (axi_spi.v/vhdl)     |         |     |
	--    |     |      |                            |         |     |
	--    |     |<---->|                            |         |     |
	--    |     |<---->|                            |         |     |
	--    |     |<---->|AXI_INTERFACE               |   SPI   |  S  |
	--    |     |<---->|                            |         |  P  |
	--    |     |<---->|                       MISO |<--------|  I  |
	--    | C   |<---->|                       MOSI |-------->|     |
	--    | P   |      |                       SCK  |-------->|     |
	--    | U   |      |                       CSn  |-------->|  D  |
	--    |     |      |                            |         |  E  |
	--    |     |----->|AXI_CLK                     |         |  V  |
	--    |     |----->|AXI_RESETn                  |         |     |
	--    |     |      |                            |         |     |
	--    |     |<-----|IRQ                         |         |     |
	--    |     |      |                            |         |     |
	--    |     |      +----------------------------+         |     |
	--    |     |                                             |     |
	--    +-----+                                             +-----+

    INST_SPI: entity work.En_SPI(Arq_SPI)
    generic map(
		C_AXI_DATA_WIDTH	=> C_AXI_DATA_WIDTH,
		C_AXI_ADDR_WIDTH	=> C_AXI_ADDR_WIDTH,
		FREQ_AXI_CLK		=> 100_000_000, -- AXI_CLK = 100MHz
		FREQ_SCLK     		=> 1_000_000)	-- SCLK = 1MHz
    port map(
		CSn			=> CSn,
		MOSI		=> MOSI,
		MISO		=> MISO,
		SCK			=> SCLK,
		INT			=> INT,
		WDATA     	=> WDATA,
		RDATA     	=> RDATA,
		WENA      	=> WENA,
		RENA      	=> RENA,
		RADDR     	=> RADDR,
		WADDR     	=> WADDR,
		AXI_CLK		=> AXI_ACLK,
		AXI_RESETn	=> AXI_ARESETN
    );
    
    ---------------------------------------------------------

end architecture arch_imp;